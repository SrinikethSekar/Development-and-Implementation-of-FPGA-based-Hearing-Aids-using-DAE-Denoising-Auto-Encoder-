module sine_wave_rom(
    input wire [9:0] addr,  // 10bit address (0 to 1023)
    output reg signed [7:0] data, // 8bit signed output
    input clk
);

    // 1024depth ROM storing sine wave values
    reg signed [7:0] rom [0:1023];

    initial begin
rom[0] = 8'd0;
rom[1] = 8'd1;
rom[2] = 8'd2;
rom[3] = 8'd2;
rom[4] = 8'd3;
rom[5] = 8'd4;
rom[6] = 8'd5;
rom[7] = 8'd5;
rom[8] = 8'd6;
rom[9] = 8'd7;
rom[10] = 8'd8;
rom[11] = 8'd9;
rom[12] = 8'd9;
rom[13] = 8'd10;
rom[14] = 8'd11;
rom[15] = 8'd12;
rom[16] = 8'd12;
rom[17] = 8'd13;
rom[18] = 8'd14;
rom[19] = 8'd15;
rom[20] = 8'd16;
rom[21] = 8'd16;
rom[22] = 8'd17;
rom[23] = 8'd18;
rom[24] = 8'd19;
rom[25] = 8'd19;
rom[26] = 8'd20;
rom[27] = 8'd21;
rom[28] = 8'd22;
rom[29] = 8'd22;
rom[30] = 8'd23;
rom[31] = 8'd24;
rom[32] = 8'd25;
rom[33] = 8'd26;
rom[34] = 8'd26;
rom[35] = 8'd27;
rom[36] = 8'd28;
rom[37] = 8'd29;
rom[38] = 8'd29;
rom[39] = 8'd30;
rom[40] = 8'd31;
rom[41] = 8'd32;
rom[42] = 8'd32;
rom[43] = 8'd33;
rom[44] = 8'd34;
rom[45] = 8'd35;
rom[46] = 8'd35;
rom[47] = 8'd36;
rom[48] = 8'd37;
rom[49] = 8'd38;
rom[50] = 8'd38;
rom[51] = 8'd39;
rom[52] = 8'd40;
rom[53] = 8'd41;
rom[54] = 8'd41;
rom[55] = 8'd42;
rom[56] = 8'd43;
rom[57] = 8'd44;
rom[58] = 8'd44;
rom[59] = 8'd45;
rom[60] = 8'd46;
rom[61] = 8'd46;
rom[62] = 8'd47;
rom[63] = 8'd48;
rom[64] = 8'd49;
rom[65] = 8'd49;
rom[66] = 8'd50;
rom[67] = 8'd51;
rom[68] = 8'd51;
rom[69] = 8'd52;
rom[70] = 8'd53;
rom[71] = 8'd54;
rom[72] = 8'd54;
rom[73] = 8'd55;
rom[74] = 8'd56;
rom[75] = 8'd56;
rom[76] = 8'd57;
rom[77] = 8'd58;
rom[78] = 8'd58;
rom[79] = 8'd59;
rom[80] = 8'd60;
rom[81] = 8'd61;
rom[82] = 8'd61;
rom[83] = 8'd62;
rom[84] = 8'd63;
rom[85] = 8'd63;
rom[86] = 8'd64;
rom[87] = 8'd65;
rom[88] = 8'd65;
rom[89] = 8'd66;
rom[90] = 8'd67;
rom[91] = 8'd67;
rom[92] = 8'd68;
rom[93] = 8'd69;
rom[94] = 8'd69;
rom[95] = 8'd70;
rom[96] = 8'd71;
rom[97] = 8'd71;
rom[98] = 8'd72;
rom[99] = 8'd72;
rom[100] = 8'd73;
rom[101] = 8'd74;
rom[102] = 8'd74;
rom[103] = 8'd75;
rom[104] = 8'd76;
rom[105] = 8'd76;
rom[106] = 8'd77;
rom[107] = 8'd78;
rom[108] = 8'd78;
rom[109] = 8'd79;
rom[110] = 8'd79;
rom[111] = 8'd80;
rom[112] = 8'd81;
rom[113] = 8'd81;
rom[114] = 8'd82;
rom[115] = 8'd82;
rom[116] = 8'd83;
rom[117] = 8'd84;
rom[118] = 8'd84;
rom[119] = 8'd85;
rom[120] = 8'd85;
rom[121] = 8'd86;
rom[122] = 8'd86;
rom[123] = 8'd87;
rom[124] = 8'd88;
rom[125] = 8'd88;
rom[126] = 8'd89;
rom[127] = 8'd89;
rom[128] = 8'd90;
rom[129] = 8'd90;
rom[130] = 8'd91;
rom[131] = 8'd91;
rom[132] = 8'd92;
rom[133] = 8'd93;
rom[134] = 8'd93;
rom[135] = 8'd94;
rom[136] = 8'd94;
rom[137] = 8'd95;
rom[138] = 8'd95;
rom[139] = 8'd96;
rom[140] = 8'd96;
rom[141] = 8'd97;
rom[142] = 8'd97;
rom[143] = 8'd98;
rom[144] = 8'd98;
rom[145] = 8'd99;
rom[146] = 8'd99;
rom[147] = 8'd100;
rom[148] = 8'd100;
rom[149] = 8'd101;
rom[150] = 8'd101;
rom[151] = 8'd102;
rom[152] = 8'd102;
rom[153] = 8'd102;
rom[154] = 8'd103;
rom[155] = 8'd103;
rom[156] = 8'd104;
rom[157] = 8'd104;
rom[158] = 8'd105;
rom[159] = 8'd105;
rom[160] = 8'd106;
rom[161] = 8'd106;
rom[162] = 8'd106;
rom[163] = 8'd107;
rom[164] = 8'd107;
rom[165] = 8'd108;
rom[166] = 8'd108;
rom[167] = 8'd109;
rom[168] = 8'd109;
rom[169] = 8'd109;
rom[170] = 8'd110;
rom[171] = 8'd110;
rom[172] = 8'd111;
rom[173] = 8'd111;
rom[174] = 8'd111;
rom[175] = 8'd112;
rom[176] = 8'd112;
rom[177] = 8'd112;
rom[178] = 8'd113;
rom[179] = 8'd113;
rom[180] = 8'd113;
rom[181] = 8'd114;
rom[182] = 8'd114;
rom[183] = 8'd114;
rom[184] = 8'd115;
rom[185] = 8'd115;
rom[186] = 8'd115;
rom[187] = 8'd116;
rom[188] = 8'd116;
rom[189] = 8'd116;
rom[190] = 8'd117;
rom[191] = 8'd117;
rom[192] = 8'd117;
rom[193] = 8'd118;
rom[194] = 8'd118;
rom[195] = 8'd118;
rom[196] = 8'd118;
rom[197] = 8'd119;
rom[198] = 8'd119;
rom[199] = 8'd119;
rom[200] = 8'd120;
rom[201] = 8'd120;
rom[202] = 8'd120;
rom[203] = 8'd120;
rom[204] = 8'd121;
rom[205] = 8'd121;
rom[206] = 8'd121;
rom[207] = 8'd121;
rom[208] = 8'd122;
rom[209] = 8'd122;
rom[210] = 8'd122;
rom[211] = 8'd122;
rom[212] = 8'd122;
rom[213] = 8'd123;
rom[214] = 8'd123;
rom[215] = 8'd123;
rom[216] = 8'd123;
rom[217] = 8'd123;
rom[218] = 8'd124;
rom[219] = 8'd124;
rom[220] = 8'd124;
rom[221] = 8'd124;
rom[222] = 8'd124;
rom[223] = 8'd124;
rom[224] = 8'd125;
rom[225] = 8'd125;
rom[226] = 8'd125;
rom[227] = 8'd125;
rom[228] = 8'd125;
rom[229] = 8'd125;
rom[230] = 8'd125;
rom[231] = 8'd126;
rom[232] = 8'd126;
rom[233] = 8'd126;
rom[234] = 8'd126;
rom[235] = 8'd126;
rom[236] = 8'd126;
rom[237] = 8'd126;
rom[238] = 8'd126;
rom[239] = 8'd126;
rom[240] = 8'd126;
rom[241] = 8'd126;
rom[242] = 8'd127;
rom[243] = 8'd127;
rom[244] = 8'd127;
rom[245] = 8'd127;
rom[246] = 8'd127;
rom[247] = 8'd127;
rom[248] = 8'd127;
rom[249] = 8'd127;
rom[250] = 8'd127;
rom[251] = 8'd127;
rom[252] = 8'd127;
rom[253] = 8'd127;
rom[254] = 8'd127;
rom[255] = 8'd127;
rom[256] = 8'd127;
rom[257] = 8'd127;
rom[258] = 8'd127;
rom[259] = 8'd127;
rom[260] = 8'd127;
rom[261] = 8'd127;
rom[262] = 8'd127;
rom[263] = 8'd127;
rom[264] = 8'd127;
rom[265] = 8'd127;
rom[266] = 8'd127;
rom[267] = 8'd127;
rom[268] = 8'd127;
rom[269] = 8'd127;
rom[270] = 8'd127;
rom[271] = 8'd126;
rom[272] = 8'd126;
rom[273] = 8'd126;
rom[274] = 8'd126;
rom[275] = 8'd126;
rom[276] = 8'd126;
rom[277] = 8'd126;
rom[278] = 8'd126;
rom[279] = 8'd126;
rom[280] = 8'd126;
rom[281] = 8'd126;
rom[282] = 8'd125;
rom[283] = 8'd125;
rom[284] = 8'd125;
rom[285] = 8'd125;
rom[286] = 8'd125;
rom[287] = 8'd125;
rom[288] = 8'd125;
rom[289] = 8'd124;
rom[290] = 8'd124;
rom[291] = 8'd124;
rom[292] = 8'd124;
rom[293] = 8'd124;
rom[294] = 8'd124;
rom[295] = 8'd123;
rom[296] = 8'd123;
rom[297] = 8'd123;
rom[298] = 8'd123;
rom[299] = 8'd123;
rom[300] = 8'd122;
rom[301] = 8'd122;
rom[302] = 8'd122;
rom[303] = 8'd122;
rom[304] = 8'd122;
rom[305] = 8'd121;
rom[306] = 8'd121;
rom[307] = 8'd121;
rom[308] = 8'd121;
rom[309] = 8'd120;
rom[310] = 8'd120;
rom[311] = 8'd120;
rom[312] = 8'd120;
rom[313] = 8'd119;
rom[314] = 8'd119;
rom[315] = 8'd119;
rom[316] = 8'd118;
rom[317] = 8'd118;
rom[318] = 8'd118;
rom[319] = 8'd118;
rom[320] = 8'd117;
rom[321] = 8'd117;
rom[322] = 8'd117;
rom[323] = 8'd116;
rom[324] = 8'd116;
rom[325] = 8'd116;
rom[326] = 8'd115;
rom[327] = 8'd115;
rom[328] = 8'd115;
rom[329] = 8'd114;
rom[330] = 8'd114;
rom[331] = 8'd114;
rom[332] = 8'd113;
rom[333] = 8'd113;
rom[334] = 8'd113;
rom[335] = 8'd112;
rom[336] = 8'd112;
rom[337] = 8'd112;
rom[338] = 8'd111;
rom[339] = 8'd111;
rom[340] = 8'd111;
rom[341] = 8'd110;
rom[342] = 8'd110;
rom[343] = 8'd109;
rom[344] = 8'd109;
rom[345] = 8'd109;
rom[346] = 8'd108;
rom[347] = 8'd108;
rom[348] = 8'd107;
rom[349] = 8'd107;
rom[350] = 8'd106;
rom[351] = 8'd106;
rom[352] = 8'd106;
rom[353] = 8'd105;
rom[354] = 8'd105;
rom[355] = 8'd104;
rom[356] = 8'd104;
rom[357] = 8'd103;
rom[358] = 8'd103;
rom[359] = 8'd102;
rom[360] = 8'd102;
rom[361] = 8'd102;
rom[362] = 8'd101;
rom[363] = 8'd101;
rom[364] = 8'd100;
rom[365] = 8'd100;
rom[366] = 8'd99;
rom[367] = 8'd99;
rom[368] = 8'd98;
rom[369] = 8'd98;
rom[370] = 8'd97;
rom[371] = 8'd97;
rom[372] = 8'd96;
rom[373] = 8'd96;
rom[374] = 8'd95;
rom[375] = 8'd95;
rom[376] = 8'd94;
rom[377] = 8'd94;
rom[378] = 8'd93;
rom[379] = 8'd93;
rom[380] = 8'd92;
rom[381] = 8'd91;
rom[382] = 8'd91;
rom[383] = 8'd90;
rom[384] = 8'd90;
rom[385] = 8'd89;
rom[386] = 8'd89;
rom[387] = 8'd88;
rom[388] = 8'd88;
rom[389] = 8'd87;
rom[390] = 8'd86;
rom[391] = 8'd86;
rom[392] = 8'd85;
rom[393] = 8'd85;
rom[394] = 8'd84;
rom[395] = 8'd84;
rom[396] = 8'd83;
rom[397] = 8'd82;
rom[398] = 8'd82;
rom[399] = 8'd81;
rom[400] = 8'd81;
rom[401] = 8'd80;
rom[402] = 8'd79;
rom[403] = 8'd79;
rom[404] = 8'd78;
rom[405] = 8'd78;
rom[406] = 8'd77;
rom[407] = 8'd76;
rom[408] = 8'd76;
rom[409] = 8'd75;
rom[410] = 8'd74;
rom[411] = 8'd74;
rom[412] = 8'd73;
rom[413] = 8'd72;
rom[414] = 8'd72;
rom[415] = 8'd71;
rom[416] = 8'd71;
rom[417] = 8'd70;
rom[418] = 8'd69;
rom[419] = 8'd69;
rom[420] = 8'd68;
rom[421] = 8'd67;
rom[422] = 8'd67;
rom[423] = 8'd66;
rom[424] = 8'd65;
rom[425] = 8'd65;
rom[426] = 8'd64;
rom[427] = 8'd63;
rom[428] = 8'd63;
rom[429] = 8'd62;
rom[430] = 8'd61;
rom[431] = 8'd61;
rom[432] = 8'd60;
rom[433] = 8'd59;
rom[434] = 8'd58;
rom[435] = 8'd58;
rom[436] = 8'd57;
rom[437] = 8'd56;
rom[438] = 8'd56;
rom[439] = 8'd55;
rom[440] = 8'd54;
rom[441] = 8'd54;
rom[442] = 8'd53;
rom[443] = 8'd52;
rom[444] = 8'd51;
rom[445] = 8'd51;
rom[446] = 8'd50;
rom[447] = 8'd49;
rom[448] = 8'd49;
rom[449] = 8'd48;
rom[450] = 8'd47;
rom[451] = 8'd46;
rom[452] = 8'd46;
rom[453] = 8'd45;
rom[454] = 8'd44;
rom[455] = 8'd44;
rom[456] = 8'd43;
rom[457] = 8'd42;
rom[458] = 8'd41;
rom[459] = 8'd41;
rom[460] = 8'd40;
rom[461] = 8'd39;
rom[462] = 8'd38;
rom[463] = 8'd38;
rom[464] = 8'd37;
rom[465] = 8'd36;
rom[466] = 8'd35;
rom[467] = 8'd35;
rom[468] = 8'd34;
rom[469] = 8'd33;
rom[470] = 8'd32;
rom[471] = 8'd32;
rom[472] = 8'd31;
rom[473] = 8'd30;
rom[474] = 8'd29;
rom[475] = 8'd29;
rom[476] = 8'd28;
rom[477] = 8'd27;
rom[478] = 8'd26;
rom[479] = 8'd26;
rom[480] = 8'd25;
rom[481] = 8'd24;
rom[482] = 8'd23;
rom[483] = 8'd22;
rom[484] = 8'd22;
rom[485] = 8'd21;
rom[486] = 8'd20;
rom[487] = 8'd19;
rom[488] = 8'd19;
rom[489] = 8'd18;
rom[490] = 8'd17;
rom[491] = 8'd16;
rom[492] = 8'd16;
rom[493] = 8'd15;
rom[494] = 8'd14;
rom[495] = 8'd13;
rom[496] = 8'd12;
rom[497] = 8'd12;
rom[498] = 8'd11;
rom[499] = 8'd10;
rom[500] = 8'd9;
rom[501] = 8'd9;
rom[502] = 8'd8;
rom[503] = 8'd7;
rom[504] = 8'd6;
rom[505] = 8'd5;
rom[506] = 8'd5;
rom[507] = 8'd4;
rom[508] = 8'd3;
rom[509] = 8'd2;
rom[510] = 8'd2;
rom[511] = 8'd1;
rom[512] = 8'd0;
rom[513] =- 8'd1;
rom[514] =- 8'd2;
rom[515] =- 8'd2;
rom[516] =- 8'd3;
rom[517] =- 8'd4;
rom[518] =- 8'd5;
rom[519] =- 8'd5;
rom[520] =- 8'd6;
rom[521] =- 8'd7;
rom[522] =- 8'd8;
rom[523] =- 8'd9;
rom[524] =- 8'd9;
rom[525] =- 8'd10;
rom[526] =- 8'd11;
rom[527] =- 8'd12;
rom[528] =- 8'd12;
rom[529] =- 8'd13;
rom[530] =- 8'd14;
rom[531] =- 8'd15;
rom[532] =- 8'd16;
rom[533] =- 8'd16;
rom[534] =- 8'd17;
rom[535] =- 8'd18;
rom[536] =- 8'd19;
rom[537] =- 8'd19;
rom[538] =- 8'd20;
rom[539] =- 8'd21;
rom[540] =- 8'd22;
rom[541] =- 8'd22;
rom[542] =- 8'd23;
rom[543] =- 8'd24;
rom[544] =- 8'd25;
rom[545] =- 8'd26;
rom[546] =- 8'd26;
rom[547] =- 8'd27;
rom[548] =- 8'd28;
rom[549] =- 8'd29;
rom[550] =- 8'd29;
rom[551] =- 8'd30;
rom[552] =- 8'd31;
rom[553] =- 8'd32;
rom[554] =- 8'd32;
rom[555] =- 8'd33;
rom[556] =- 8'd34;
rom[557] =- 8'd35;
rom[558] =- 8'd35;
rom[559] =- 8'd36;
rom[560] =- 8'd37;
rom[561] =- 8'd38;
rom[562] =- 8'd38;
rom[563] =- 8'd39;
rom[564] =- 8'd40;
rom[565] =- 8'd41;
rom[566] =- 8'd41;
rom[567] =- 8'd42;
rom[568] =- 8'd43;
rom[569] =- 8'd44;
rom[570] =- 8'd44;
rom[571] =- 8'd45;
rom[572] =- 8'd46;
rom[573] =- 8'd46;
rom[574] =- 8'd47;
rom[575] =- 8'd48;
rom[576] =- 8'd49;
rom[577] =- 8'd49;
rom[578] =- 8'd50;
rom[579] =- 8'd51;
rom[580] =- 8'd51;
rom[581] =- 8'd52;
rom[582] =- 8'd53;
rom[583] =- 8'd54;
rom[584] =- 8'd54;
rom[585] =- 8'd55;
rom[586] =- 8'd56;
rom[587] =- 8'd56;
rom[588] =- 8'd57;
rom[589] =- 8'd58;
rom[590] =- 8'd58;
rom[591] =- 8'd59;
rom[592] =- 8'd60;
rom[593] =- 8'd61;
rom[594] =- 8'd61;
rom[595] =- 8'd62;
rom[596] =- 8'd63;
rom[597] =- 8'd63;
rom[598] =- 8'd64;
rom[599] =- 8'd65;
rom[600] =- 8'd65;
rom[601] =- 8'd66;
rom[602] =- 8'd67;
rom[603] =- 8'd67;
rom[604] =- 8'd68;
rom[605] =- 8'd69;
rom[606] =- 8'd69;
rom[607] =- 8'd70;
rom[608] =- 8'd71;
rom[609] =- 8'd71;
rom[610] =- 8'd72;
rom[611] =- 8'd72;
rom[612] =- 8'd73;
rom[613] =- 8'd74;
rom[614] =- 8'd74;
rom[615] =- 8'd75;
rom[616] =- 8'd76;
rom[617] =- 8'd76;
rom[618] =- 8'd77;
rom[619] =- 8'd78;
rom[620] =- 8'd78;
rom[621] =- 8'd79;
rom[622] =- 8'd79;
rom[623] =- 8'd80;
rom[624] =- 8'd81;
rom[625] =- 8'd81;
rom[626] =- 8'd82;
rom[627] =- 8'd82;
rom[628] =- 8'd83;
rom[629] =- 8'd84;
rom[630] =- 8'd84;
rom[631] =- 8'd85;
rom[632] =- 8'd85;
rom[633] =- 8'd86;
rom[634] =- 8'd86;
rom[635] =- 8'd87;
rom[636] =- 8'd88;
rom[637] =- 8'd88;
rom[638] =- 8'd89;
rom[639] =- 8'd89;
rom[640] =- 8'd90;
rom[641] =- 8'd90;
rom[642] =- 8'd91;
rom[643] =- 8'd91;
rom[644] =- 8'd92;
rom[645] =- 8'd93;
rom[646] =- 8'd93;
rom[647] =- 8'd94;
rom[648] =- 8'd94;
rom[649] =- 8'd95;
rom[650] =- 8'd95;
rom[651] =- 8'd96;
rom[652] =- 8'd96;
rom[653] =- 8'd97;
rom[654] =- 8'd97;
rom[655] =- 8'd98;
rom[656] =- 8'd98;
rom[657] =- 8'd99;
rom[658] =- 8'd99;
rom[659] =- 8'd100;
rom[660] =- 8'd100;
rom[661] =- 8'd101;
rom[662] =- 8'd101;
rom[663] =- 8'd102;
rom[664] =- 8'd102;
rom[665] =- 8'd102;
rom[666] =- 8'd103;
rom[667] =- 8'd103;
rom[668] =- 8'd104;
rom[669] =- 8'd104;
rom[670] =- 8'd105;
rom[671] =- 8'd105;
rom[672] =- 8'd106;
rom[673] =- 8'd106;
rom[674] =- 8'd106;
rom[675] =- 8'd107;
rom[676] =- 8'd107;
rom[677] =- 8'd108;
rom[678] =- 8'd108;
rom[679] =- 8'd109;
rom[680] =- 8'd109;
rom[681] =- 8'd109;
rom[682] =- 8'd110;
rom[683] =- 8'd110;
rom[684] =- 8'd111;
rom[685] =- 8'd111;
rom[686] =- 8'd111;
rom[687] =- 8'd112;
rom[688] =- 8'd112;
rom[689] =- 8'd112;
rom[690] =- 8'd113;
rom[691] =- 8'd113;
rom[692] =- 8'd113;
rom[693] =- 8'd114;
rom[694] =- 8'd114;
rom[695] =- 8'd114;
rom[696] =- 8'd115;
rom[697] =- 8'd115;
rom[698] =- 8'd115;
rom[699] =- 8'd116;
rom[700] =- 8'd116;
rom[701] =- 8'd116;
rom[702] =- 8'd117;
rom[703] =- 8'd117;
rom[704] =- 8'd117;
rom[705] =- 8'd118;
rom[706] =- 8'd118;
rom[707] =- 8'd118;
rom[708] =- 8'd118;
rom[709] =- 8'd119;
rom[710] =- 8'd119;
rom[711] =- 8'd119;
rom[712] =- 8'd120;
rom[713] =- 8'd120;
rom[714] =- 8'd120;
rom[715] =- 8'd120;
rom[716] =- 8'd121;
rom[717] =- 8'd121;
rom[718] =- 8'd121;
rom[719] =- 8'd121;
rom[720] =- 8'd122;
rom[721] =- 8'd122;
rom[722] =- 8'd122;
rom[723] =- 8'd122;
rom[724] =- 8'd122;
rom[725] =- 8'd123;
rom[726] =- 8'd123;
rom[727] =- 8'd123;
rom[728] =- 8'd123;
rom[729] =- 8'd123;
rom[730] =- 8'd124;
rom[731] =- 8'd124;
rom[732] =- 8'd124;
rom[733] =- 8'd124;
rom[734] =- 8'd124;
rom[735] =- 8'd124;
rom[736] =- 8'd125;
rom[737] =- 8'd125;
rom[738] =- 8'd125;
rom[739] =- 8'd125;
rom[740] =- 8'd125;
rom[741] =- 8'd125;
rom[742] =- 8'd125;
rom[743] =- 8'd126;
rom[744] =- 8'd126;
rom[745] =- 8'd126;
rom[746] =- 8'd126;
rom[747] =- 8'd126;
rom[748] =- 8'd126;
rom[749] =- 8'd126;
rom[750] =- 8'd126;
rom[751] =- 8'd126;
rom[752] =- 8'd126;
rom[753] =- 8'd126;
rom[754] =- 8'd127;
rom[755] =- 8'd127;
rom[756] =- 8'd127;
rom[757] =- 8'd127;
rom[758] =- 8'd127;
rom[759] =- 8'd127;
rom[760] =- 8'd127;
rom[761] =- 8'd127;
rom[762] =- 8'd127;
rom[763] =- 8'd127;
rom[764] =- 8'd127;
rom[765] =- 8'd127;
rom[766] =- 8'd127;
rom[767] =- 8'd127;
rom[768] =- 8'd127;
rom[769] =- 8'd127;
rom[770] =- 8'd127;
rom[771] =- 8'd127;
rom[772] =- 8'd127;
rom[773] =- 8'd127;
rom[774] =- 8'd127;
rom[775] =- 8'd127;
rom[776] =- 8'd127;
rom[777] =- 8'd127;
rom[778] =- 8'd127;
rom[779] =- 8'd127;
rom[780] =- 8'd127;
rom[781] =- 8'd127;
rom[782] =- 8'd127;
rom[783] =- 8'd126;
rom[784] =- 8'd126;
rom[785] =- 8'd126;
rom[786] =- 8'd126;
rom[787] =- 8'd126;
rom[788] =- 8'd126;
rom[789] =- 8'd126;
rom[790] =- 8'd126;
rom[791] =- 8'd126;
rom[792] =- 8'd126;
rom[793] =- 8'd126;
rom[794] =- 8'd125;
rom[795] =- 8'd125;
rom[796] =- 8'd125;
rom[797] =- 8'd125;
rom[798] =- 8'd125;
rom[799] =- 8'd125;
rom[800] =- 8'd125;
rom[801] =- 8'd124;
rom[802] =- 8'd124;
rom[803] =- 8'd124;
rom[804] =- 8'd124;
rom[805] =- 8'd124;
rom[806] =- 8'd124;
rom[807] =- 8'd123;
rom[808] =- 8'd123;
rom[809] =- 8'd123;
rom[810] =- 8'd123;
rom[811] =- 8'd123;
rom[812] =- 8'd122;
rom[813] =- 8'd122;
rom[814] =- 8'd122;
rom[815] =- 8'd122;
rom[816] =- 8'd122;
rom[817] =- 8'd121;
rom[818] =- 8'd121;
rom[819] =- 8'd121;
rom[820] =- 8'd121;
rom[821] =- 8'd120;
rom[822] =- 8'd120;
rom[823] =- 8'd120;
rom[824] =- 8'd120;
rom[825] =- 8'd119;
rom[826] =- 8'd119;
rom[827] =- 8'd119;
rom[828] =- 8'd118;
rom[829] =- 8'd118;
rom[830] =- 8'd118;
rom[831] =- 8'd118;
rom[832] =- 8'd117;
rom[833] =- 8'd117;
rom[834] =- 8'd117;
rom[835] =- 8'd116;
rom[836] =- 8'd116;
rom[837] =- 8'd116;
rom[838] =- 8'd115;
rom[839] =- 8'd115;
rom[840] =- 8'd115;
rom[841] =- 8'd114;
rom[842] =- 8'd114;
rom[843] =- 8'd114;
rom[844] =- 8'd113;
rom[845] =- 8'd113;
rom[846] =- 8'd113;
rom[847] =- 8'd112;
rom[848] =- 8'd112;
rom[849] =- 8'd112;
rom[850] =- 8'd111;
rom[851] =- 8'd111;
rom[852] =- 8'd111;
rom[853] =- 8'd110;
rom[854] =- 8'd110;
rom[855] =- 8'd109;
rom[856] =- 8'd109;
rom[857] =- 8'd109;
rom[858] =- 8'd108;
rom[859] =- 8'd108;
rom[860] =- 8'd107;
rom[861] =- 8'd107;
rom[862] =- 8'd106;
rom[863] =- 8'd106;
rom[864] =- 8'd106;
rom[865] =- 8'd105;
rom[866] =- 8'd105;
rom[867] =- 8'd104;
rom[868] =- 8'd104;
rom[869] =- 8'd103;
rom[870] =- 8'd103;
rom[871] =- 8'd102;
rom[872] =- 8'd102;
rom[873] =- 8'd102;
rom[874] =- 8'd101;
rom[875] =- 8'd101;
rom[876] =- 8'd100;
rom[877] =- 8'd100;
rom[878] =- 8'd99;
rom[879] =- 8'd99;
rom[880] =- 8'd98;
rom[881] =- 8'd98;
rom[882] =- 8'd97;
rom[883] =- 8'd97;
rom[884] =- 8'd96;
rom[885] =- 8'd96;
rom[886] =- 8'd95;
rom[887] =- 8'd95;
rom[888] =- 8'd94;
rom[889] =- 8'd94;
rom[890] =- 8'd93;
rom[891] =- 8'd93;
rom[892] =- 8'd92;
rom[893] =- 8'd91;
rom[894] =- 8'd91;
rom[895] =- 8'd90;
rom[896] =- 8'd90;
rom[897] =- 8'd89;
rom[898] =- 8'd89;
rom[899] =- 8'd88;
rom[900] =- 8'd88;
rom[901] =- 8'd87;
rom[902] =- 8'd86;
rom[903] =- 8'd86;
rom[904] =- 8'd85;
rom[905] =- 8'd85;
rom[906] =- 8'd84;
rom[907] =- 8'd84;
rom[908] =- 8'd83;
rom[909] =- 8'd82;
rom[910] =- 8'd82;
rom[911] =- 8'd81;
rom[912] =- 8'd81;
rom[913] =- 8'd80;
rom[914] =- 8'd79;
rom[915] =- 8'd79;
rom[916] =- 8'd78;
rom[917] =- 8'd78;
rom[918] =- 8'd77;
rom[919] =- 8'd76;
rom[920] =- 8'd76;
rom[921] =- 8'd75;
rom[922] =- 8'd74;
rom[923] =- 8'd74;
rom[924] =- 8'd73;
rom[925] =- 8'd72;
rom[926] =- 8'd72;
rom[927] =- 8'd71;
rom[928] =- 8'd71;
rom[929] =- 8'd70;
rom[930] =- 8'd69;
rom[931] =- 8'd69;
rom[932] =- 8'd68;
rom[933] =- 8'd67;
rom[934] =- 8'd67;
rom[935] =- 8'd66;
rom[936] =- 8'd65;
rom[937] =- 8'd65;
rom[938] =- 8'd64;
rom[939] =- 8'd63;
rom[940] =- 8'd63;
rom[941] =- 8'd62;
rom[942] =- 8'd61;
rom[943] =- 8'd61;
rom[944] =- 8'd60;
rom[945] =- 8'd59;
rom[946] =- 8'd58;
rom[947] =- 8'd58;
rom[948] =- 8'd57;
rom[949] =- 8'd56;
rom[950] =- 8'd56;
rom[951] =- 8'd55;
rom[952] =- 8'd54;
rom[953] =- 8'd54;
rom[954] =- 8'd53;
rom[955] =- 8'd52;
rom[956] =- 8'd51;
rom[957] =- 8'd51;
rom[958] =- 8'd50;
rom[959] =- 8'd49;
rom[960] =- 8'd49;
rom[961] =- 8'd48;
rom[962] =- 8'd47;
rom[963] =- 8'd46;
rom[964] =- 8'd46;
rom[965] =- 8'd45;
rom[966] =- 8'd44;
rom[967] =- 8'd44;
rom[968] =- 8'd43;
rom[969] =- 8'd42;
rom[970] =- 8'd41;
rom[971] =- 8'd41;
rom[972] =- 8'd40;
rom[973] =- 8'd39;
rom[974] =- 8'd38;
rom[975] =- 8'd38;
rom[976] =- 8'd37;
rom[977] =- 8'd36;
rom[978] =- 8'd35;
rom[979] =- 8'd35;
rom[980] =- 8'd34;
rom[981] =- 8'd33;
rom[982] =- 8'd32;
rom[983] =- 8'd32;
rom[984] =- 8'd31;
rom[985] =- 8'd30;
rom[986] =- 8'd29;
rom[987] =- 8'd29;
rom[988] =- 8'd28;
rom[989] =- 8'd27;
rom[990] =- 8'd26;
rom[991] =- 8'd26;
rom[992] =- 8'd25;
rom[993] =- 8'd24;
rom[994] =- 8'd23;
rom[995] =- 8'd22;
rom[996] =- 8'd22;
rom[997] =- 8'd21;
rom[998] =- 8'd20;
rom[999] =- 8'd19;
rom[1000] =- 8'd19;
rom[1001] =- 8'd18;
rom[1002] =- 8'd17;
rom[1003] =- 8'd16;
rom[1004] =- 8'd16;
rom[1005] =- 8'd15;
rom[1006] =- 8'd14;
rom[1007] =- 8'd13;
rom[1008] =- 8'd12;
rom[1009] =- 8'd12;
rom[1010] =- 8'd11;
rom[1011] =- 8'd10;
rom[1012] =- 8'd9;
rom[1013] =- 8'd9;
rom[1014] =- 8'd8;
rom[1015] =- 8'd7;
rom[1016] =- 8'd6;
rom[1017] =- 8'd5;
rom[1018] =- 8'd5;
rom[1019] =- 8'd4;
rom[1020] =- 8'd3;
rom[1021] =- 8'd2;
rom[1022] =- 8'd2;
rom[1023] =- 8'd1;
 end

    always @(clk) begin
        data = rom[addr];
    end

endmodule
